module small_pseudo_cpu